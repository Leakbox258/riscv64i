module top (
    input i_clk,
    input i_rst,
    output [15:0] o_ledr,
);


endmodule