`include "pipeline_pkg.sv"

module ControlFlowPredict
  import pipeline_pkg::*;
();

endmodule
