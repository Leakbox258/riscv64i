module MEM #(
    DATA_WIDTH = 64
) ();

endmodule
